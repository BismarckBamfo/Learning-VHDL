----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:33:16 01/22/2020 
-- Design Name: 
-- Module Name:    sys1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sys1 is
    Port ( a_in1 : in  STD_LOGIC;
           b_in2 : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           ctrl_int : in  STD_LOGIC;
           out_b : out  STD_LOGIC);
end sys1;

architecture Behavioral of sys1 is

begin


end Behavioral;

