----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:05:00 02/14/2020 
-- Design Name: 
-- Module Name:    my_ckt - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity my_ckt is
	port (
				A,B,c : IN STD_LOGIC;
				Y		: OUT STD_LOGIC
			);
end my_ckt;

architecture Behavioral of my_ckt is

begin
	my_ckt : process(b) 
					begin 
						Y <= (A and B ) OR (A nand C);
					end process;
	

end Behavioral;

