----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:10:46 02/26/2020 
-- Design Name: 
-- Module Name:    case_Mux_8to1_testcase - case_Mux_8to1_testcase_OP 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity case_Mux_8to1_testcase is
end case_Mux_8to1_testcase;

architecture case_Mux_8to1_testcase_OP of case_Mux_8to1_testcase is

begin


end case_Mux_8to1_testcase_OP;

